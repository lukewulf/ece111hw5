import definitions::*;

module FPU_D();

endmodule
